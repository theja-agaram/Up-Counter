* C:\Users\theja\Desktop\counter.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/04/22 00:05:07

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  ? ? ? ? ? Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ ? ? ? ? theja_async4bitupcounter		
U8  Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_R6-Pad1_ O1 O2 O3 dac_bridge_4		
U7  clock rst3 rst2 ? rst0 ? ? ? ? ? adc_bridge_5		
R6  Net-_R6-Pad1_ Net-_C1-Pad1_ 1k		
R2  Net-_R2-Pad1_ clock 1k		
R1  Net-_R1-Pad1_ rst3 1k		
R3  rst2 Net-_R3-Pad2_ 1k		
R4  rst1 Net-_R4-Pad2_ 1k		
R5  rst0 Net-_R5-Pad2_ 1k		
C1  Net-_C1-Pad1_ GND 1u		
v1  Net-_R2-Pad1_ GND pulse		
v2  Net-_R1-Pad1_ GND pulse		
v3  Net-_R3-Pad2_ GND pulse		
v4  Net-_R4-Pad2_ GND pulse		
v5  Net-_R5-Pad2_ GND pulse		
U9  Net-_C1-Pad1_ plot_v1		
U10  O1 plot_v1		
U11  O2 plot_v1		
U12  O3 plot_v1		
U2  clock plot_v1		
U3  rst3 plot_v1		
U4  rst2 plot_v1		
U5  rst1 plot_v1		
U6  rst0 plot_v1		

.end
